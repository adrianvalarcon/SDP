----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01/29/2021 02:39:46 AM
-- Design Name: 
-- Module Name: uart_rx - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity uart_rx is
    generic (
        D_bit   : integer := 8;     -- # of data bits
        SB_tick : integer := 16     -- # of ticks for stop bits (2 * # stop bits)
    );
    
    port (
        clk     : in  std_logic;
        reset   : in  std_logic;
        rx      : in  std_logic;                    -- Receive data bit
        s_tick  : in  std_logic;                    -- Start flag
        rx_done : out std_logic;                    -- Done flag
        d_out   : out std_logic_vector(7 downto 0)  -- 8 data bits
    );
end uart_rx;

architecture Behavioral of uart_rx is
    type state_type is (idle, start, data, stop);
    signal state_reg, state_next : state_type;
    signal s_reg, s_next : unsigned(3 downto 0);        -- State registers
    signal n_reg, n_next : unsigned(2 downto 0);        -- Data bit position register
    signal b_reg, b_next : std_logic_vector(7 downto 0);-- 

begin
    
    -- FSMD state/data regs
    process(clk, reset)
    begin
        if (reset = '1') then
            state_reg <= idle;
            s_reg <= (others => '0');
            n_reg <= (others => '0');
            b_reg <= (others => '0');
        elsif (clk'event and clk = '1') then
            state_reg <= state_next;
            s_reg <= s_next;
            n_reg <= n_next;
            b_reg <= b_next;
        end if;
    end process;

    -- Next state logic
    process (state_reg, s_reg, n_reg, b_reg, s_tick, rx)
    begin
        state_next  <= state_reg;
        s_next      <= s_reg;
        n_next      <= n_reg;
        b_next      <= b_reg;
        rx_done     <= '0';
        
        case state_reg is
            -- Idle state
            when idle =>
                if (rx = '0') then
                    state_next <= start;
                    s_next <= (others => '0');
                end if;
            
            -- Start receive sequence
            when start =>
                if (s_tick = '1') then
                    if (s_reg = 7) then
                        state_next <= data;
                        s_next <= (others => '0');
                        n_next <= (others => '0');
                    else
                        s_next <= s_reg + 1;
                    end if;
                end if;
                
            -- Receive Data
            when data =>
                if (s_tick = '1') then
                    if (s_reg = 15) then
                        s_next <= (others => '0');
                        b_next <= rx & b_reg(7 downto 1);
                        if (n_reg = (D_bit - 1)) then
                            state_next <= stop;
                        else
                            n_next <= n_reg + 1;
                        end if;
                    else
                        s_next <= s_reg + 1;
                    end if;
                end if;
                    
            -- Stop receiving
            when stop =>
                if (s_tick = '1') then
                    if (s_reg = (SB_tick - 1)) then
                        state_next <= idle;
                        rx_done <= '1';
                    else
                        s_next <= s_reg + 1;
                    end if;
                end if;
                
        end case;
    end process;
    
    -- Output received data bits
    d_out <= b_reg;
    
end Behavioral;